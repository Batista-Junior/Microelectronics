CIRCUIT C:\Users\Batista\Desktop\MEU_TRABALHO_FINAL\OSCILATOR_RING\OSC_RING_7.MSK
*
* IC Technology: CMOS 90nm, 6 Metal Copper - strained SiGe - LowK
*
VDD 1 0 DC 1.20
*
* List of nodes
* "S_1" corresponds to n�3
* "S_7" corresponds to n�5
* "S_6" corresponds to n�6
* "S_5" corresponds to n�7
* "S_4" corresponds to n�8
* "S_3" corresponds to n�9
* "S_2" corresponds to n�10
*
* MOS devices
MN1 0 5 3 0 N1  W= 0.60U L= 0.10U
MN2 0 6 5 0 N1  W= 0.60U L= 0.10U
MN3 0 7 6 0 N1  W= 0.60U L= 0.10U
MN4 0 8 7 0 N1  W= 0.60U L= 0.10U
MN5 0 9 8 0 N1  W= 0.60U L= 0.10U
MN6 0 10 9 0 N1  W= 0.60U L= 0.10U
MN7 0 3 10 0 N1  W= 0.60U L= 0.10U
MP1 1 5 3 1 P1  W= 1.00U L= 0.10U
MP2 1 6 5 1 P1  W= 1.00U L= 0.10U
MP3 1 7 6 1 P1  W= 1.00U L= 0.10U
MP4 1 8 7 1 P1  W= 1.00U L= 0.10U
MP5 1 9 8 1 P1  W= 1.00U L= 0.10U
MP6 1 10 9 1 P1  W= 1.00U L= 0.10U
MP7 1 3 10 1 P1  W= 1.00U L= 0.10U
*
C2 1 0  2.400fF
C3 3 0  1.205fF
C4 1 0  3.013fF
C5 5 0  0.646fF
C6 6 0  0.646fF
C7 7 0  0.646fF
C8 8 0  0.646fF
C9 9 0  0.629fF
C10 10 0  0.629fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.28 U0=0.060 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  0.9 U0=0.060 UA=3.400e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.32 U0=0.027 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.9 U0=0.027 UA=2.200e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 2.00N
print  V(3) V(10) V(9) V(8) V(7) V(6) V(5) > out.txt
plot  V(3) V(10) V(9) V(8) V(7) V(6) V(5)
.endc
.END
