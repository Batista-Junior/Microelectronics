CIRCUIT C:\Users\Batista\Desktop\RESIDENCIA_EM_MICROELETRONICA\MICROWIND\TRINAND\TRINAND_MWIND.MSK
*
* IC Technology: CMOS 90nm, 6 Metal Copper - strained SiGe - LowK
*
VDD 1 0 DC 1.20
VC 8 0 DC 0 PULSE(0.00 1.20 0.79N 0.01N 0.01N 0.79N 1.60N)
VA 9 0 DC 0 PULSE(0.00 1.20 0.17N 0.01N 0.01N 0.17N 0.36N)
VB 10 0 DC 0 PULSE(0.00 1.20 0.39N 0.01N 0.01N 0.39N 0.80N)
*
* List of nodes
* "Y" corresponds to n�3
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "C" corresponds to n�8
* "A" corresponds to n�9
* "B" corresponds to n�10
*
* MOS devices
MN1 5 8 3 0 N1  W= 0.60U L= 0.10U
MN2 6 10 5 0 N1  W= 0.60U L= 0.10U
MN3 0 9 6 0 N1  W= 0.60U L= 0.10U
MP1 1 8 3 1 P1  W= 0.60U L= 0.10U
MP2 3 10 1 1 P1  W= 0.60U L= 0.10U
MP3 1 9 3 1 P1  W= 0.60U L= 0.10U
*
C2 1 0  0.600fF
C3 3 0  0.868fF
C4 1 0  0.611fF
C5 5 0  0.153fF
C6 6 0  0.153fF
C8 8 0  0.058fF
C9 9 0  0.058fF
C10 10 0  0.058fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.28 U0=0.060 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  0.9 U0=0.060 UA=3.400e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.32 U0=0.027 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.9 U0=0.027 UA=2.200e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 5.00N
print  V(8) V(3) V(9) V(10) > out.txt
plot  V(8) V(3) V(9) V(10)
.endc
.END
